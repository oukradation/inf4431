library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
entity p_ctrl is
  port (
    -- System Clock and Reset
    rst_div       : in  std_logic;           -- Reset
    mclk_div       : in  std_logic;           -- Clock
    sp        : in  signed(7 downto 0);  -- Set Point
    pos       : in  signed(7 downto 0);  -- Measured position
    motor_cw  : out std_logic;           --Motor Clock Wise direction
    motor_ccw : out std_logic            --Motor Counter Clock Wise direction
    );      
end entity;
